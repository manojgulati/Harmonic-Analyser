-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Sunday, November 16, 2014 00:40:24 India Standard Time

